localparam PTR_RESET = 0;
localparam PTR_PAUSE = 1;
localparam PTR_START = 2;
localparam PTR_RIGHT = 4;
localparam PTR_LEFT = 5;

localparam MEM_WRITE = 0;
localparam MEM_READ = 1;
localparam MEM_ECHO = 2;
