localparam PTR_RESET = 0
localparam PTR_PAUSE = 1;
localparam PTR_START = 2;
localparam PTR_RIGHT = 3;
localparam PTR_LEFT = 4;

localparam MEM_WRITE = 0;
localparam MEM_READ = 1;
