localparam PTR_PAUSE = 0;
localparam PTR_START = 1;
localparam PTR_RESET = 2;

localparam MEM_WRITE = 0;
localparam MEM_READ = 1;
